module top_module(
    input clk,
    input load,
    input [1:0] ena,
    input [99:0] data,
    output reg [99:0] q); 
    
    parameter N = 99;   // number of bits - 1  // for scalable code
    always @(posedge clk)begin
        if (load) q <= data;
        else case(ena)
            2'b01: q <= {q[0], q[N:1]};
            2'b10: q <= {q[N-1:0],q[N]};
        endcase
    end

endmodule
