module top_module (
    input clk,
    input resetn,
    input [1:0] byteena,
    input [15:0] d,
    output [15:0] q
);
    always @(posedge clk)
        if (!resetn) q <= 16'b0;
    	else begin 
            q[7:0] <= byteena[0] ? d[7:0] : q[7:0];
            q[15:8] <= byteena[1] ? d[15:8] : q[15:8];
        end
  
//  since we are intentionally creating flip flops hence we shall not else logic 
  // m = 2: 
  /*
      always @(posedge clk)
        begin
            if (!resetn) q <= 16'b0 ;
            else begin
                if (byteena[1]) q[15:8] <= d[15:8];
                if (byteena[0]) q[7:0] <= d[7:0];
            end
    */

endmodule
